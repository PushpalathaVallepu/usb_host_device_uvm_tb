`ifndef USB_HOST_XFER_ITEM_SV
  `define USB_HOST_XFER_ITEM_SV

typedef enum {USB_SOF, USB_OUT, USB_IN, USB_SETUP, ACK} usb_xfer_type_e;

class usb_host_xfer_item extends uvm_sequence_item;

  usb_xfer_type_e xfer_type;

  // Packet handles
  rand sof_pkt    sof;
  rand token_pkt  token;
  rand data_pkt   data;
  rand hs_pkt     hs;

  // Queues for coverage or test expansion
  rand token_pkt  tokenQ[$];
  rand data_pkt   dataQ[$];
  rand hs_pkt     hsQ[$];

  // I/O helper fields
  bit [7:0] dout;
  bit [7:0] din;

  // Serialized byte stream
  byte unsigned tx_bytes[$];
  byte unsigned rx_bytes[$];

  // ----------------------------------------------------------
  // Factory registration
  // ----------------------------------------------------------
  `uvm_object_utils_begin(usb_host_xfer_item)
    `uvm_field_enum        (usb_xfer_type_e, xfer_type, UVM_DEFAULT)
    `uvm_field_object      (sof,      UVM_DEFAULT)
    `uvm_field_object      (token,    UVM_DEFAULT)
    `uvm_field_object      (data,     UVM_DEFAULT)
    `uvm_field_object      (hs,       UVM_DEFAULT)
    `uvm_field_queue_object(tokenQ,   UVM_DEFAULT)
    `uvm_field_queue_object(dataQ,    UVM_DEFAULT)
    `uvm_field_queue_object(hsQ,      UVM_DEFAULT)
  `uvm_object_utils_end

  // ----------------------------------------------------------
  function new(string name = "usb_host_xfer_item");
    super.new(name);
  endfunction

  // ----------------------------------------------------------
  function void pre_randomize();
    sof   = sof_pkt   ::type_id::create("sof");
    token = token_pkt ::type_id::create("token");
    data  = data_pkt  ::type_id::create("data");
    hs    = hs_pkt    ::type_id::create("hs");

    tokenQ.delete();
    dataQ.delete();
    hsQ.delete();

    tokenQ.push_back(token_pkt::type_id::create("tokenQ[0]"));
    dataQ.push_back(data_pkt ::type_id::create("dataQ[0]"));
    hsQ  .push_back(hs_pkt   ::type_id::create("hsQ[0]"));
  endfunction

  // ----------------------------------------------------------
  function void post_randomize();
    xfer_type = usb_decode_pid(token.pid);
  endfunction

  // ----------------------------------------------------------
function string convert2string();
  string s;
  s = $sformatf("xfer_type=%s | ", xfer_type.name());

  if (tokenQ.size() > 0)
    s = {s, $sformatf("token: pid=0x%0h addr=%0d ep=%0d | ",
        token.pid, token.addr, token.ep_no)};
  else
    s = {s, "token: N/A | "};

  case (xfer_type)
    USB_OUT, USB_SETUP: begin
      if (dataQ.size() > 0)
        s = {s, $sformatf("data: pid=0x%0h len=%0d | ",
          data.pid, data.dataQ.size())};
      else
        s = {s, "data: N/A | "};

      if (hsQ.size() > 0)
        s = {s, $sformatf("handshake: pid=0x%0h", hs.pid)};
      else
        s = {s, "handshake: N/A"};
    end

    USB_IN: begin
      if (hsQ.size() > 0)
        s = {s, $sformatf("handshake: pid=0x%0h | ", hs.pid)};
      else
        s = {s, "handshake: N/A | "};

      if (dataQ.size() > 0)
        s = {s, $sformatf("data: pid=0x%0h len=%0d",
          data.pid, data.dataQ.size())};
      else
        s = {s, "data: N/A"};
    end

    USB_SOF: begin
      s = {s, "Start-of-Frame only"};
    end

    default: s = {s, "Unknown transfer"};
  endcase

  return s;
endfunction
  
  //------------------------------------------------------------------
  // serialise host generated bytes into tx_bytes[$]
  //------------------------------------------------------------------
function void pack_for_host();
  tx_bytes.delete();

  case (xfer_type)
    USB_SOF: begin
      tx_bytes.push_back(sof.pid);                        // PID
      tx_bytes.push_back(sof.frame_no[7:0]);              // Frame number LSB
      tx_bytes.push_back({sof.crc, sof.frame_no[10:8]});  // CRC5 + upper frame bits
    end

    USB_OUT, USB_SETUP: begin
      tx_bytes.push_back(token.pid);                             // PID
      tx_bytes.push_back({token.addr});                          // Address (7 bits)
      tx_bytes.push_back({token.crc, token.ep_no[3:1]});         // CRC5 + upper EP bits
      tx_bytes.push_back(data.pid);                              // DATA PID
      foreach (data.dataQ[i]) tx_bytes.push_back(data.dataQ[i]); // Payload
      tx_bytes.push_back(data.crc[7:0]);                         // CRC16 LSB
      tx_bytes.push_back(data.crc[15:8]);                        // CRC16 MSB
    end

    USB_IN: begin
      tx_bytes.push_back(token.pid);                             // PID
      tx_bytes.push_back({token.addr});                          // Address
      tx_bytes.push_back({token.crc, token.ep_no[3:1]});         // CRC5 + EP
      // IN: Expect response from device later
    end

    default: begin
      `uvm_warning("PACK", "Unknown transfer type in pack_for_host()")
    end
  endcase
endfunction
function automatic usb_xfer_type_e usb_decode_pid(byte pid);
  case (pid[3:0]) // lower 4 bits
    4'h1: return USB_OUT;
    4'h9: return USB_IN;
    4'hD: return USB_SETUP;
    4'h5: return USB_SOF;
    4'h2: return ACK;
    default: $display("UNKNOWN");
  endcase
endfunction
  
endclass

`endif
